module aes_sbox_v3 (dec,
    S,
    U);
 input dec;
 output [7:0] S;
 input [7:0] U;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;

 sky130_fd_sc_hd__buf_4 _262_ (.A(net4),
    .X(_089_));
 sky130_fd_sc_hd__clkbuf_4 _263_ (.A(net2),
    .X(_100_));
 sky130_fd_sc_hd__xnor2_4 _264_ (.A(_089_),
    .B(_100_),
    .Y(_111_));
 sky130_fd_sc_hd__buf_4 _265_ (.A(net7),
    .X(_121_));
 sky130_fd_sc_hd__xor2_4 _266_ (.A(_121_),
    .B(net6),
    .X(_132_));
 sky130_fd_sc_hd__xor2_1 _267_ (.A(_111_),
    .B(_132_),
    .X(_142_));
 sky130_fd_sc_hd__xnor2_4 _268_ (.A(net3),
    .B(net6),
    .Y(_152_));
 sky130_fd_sc_hd__xor2_1 _269_ (.A(_111_),
    .B(_152_),
    .X(_162_));
 sky130_fd_sc_hd__clkinv_2 _270_ (.A(net9),
    .Y(_172_));
 sky130_fd_sc_hd__mux2_1 _271_ (.A0(_142_),
    .A1(_162_),
    .S(_172_),
    .X(_182_));
 sky130_fd_sc_hd__buf_2 _272_ (.A(net9),
    .X(_190_));
 sky130_fd_sc_hd__buf_2 _273_ (.A(_190_),
    .X(_191_));
 sky130_fd_sc_hd__buf_6 _274_ (.A(net5),
    .X(_192_));
 sky130_fd_sc_hd__xnor2_4 _275_ (.A(_192_),
    .B(_089_),
    .Y(_193_));
 sky130_fd_sc_hd__clkbuf_4 _276_ (.A(net8),
    .X(_194_));
 sky130_fd_sc_hd__xor2_4 _277_ (.A(_192_),
    .B(_194_),
    .X(_195_));
 sky130_fd_sc_hd__nor2_1 _278_ (.A(_190_),
    .B(_195_),
    .Y(_196_));
 sky130_fd_sc_hd__a21oi_2 _279_ (.A1(_191_),
    .A2(_193_),
    .B1(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__clkbuf_4 _280_ (.A(_172_),
    .X(_198_));
 sky130_fd_sc_hd__xor2_1 _281_ (.A(net3),
    .B(_100_),
    .X(_199_));
 sky130_fd_sc_hd__xnor2_1 _282_ (.A(_193_),
    .B(_199_),
    .Y(_200_));
 sky130_fd_sc_hd__xor2_2 _283_ (.A(_194_),
    .B(_121_),
    .X(_201_));
 sky130_fd_sc_hd__buf_4 _284_ (.A(net1),
    .X(_202_));
 sky130_fd_sc_hd__xor2_2 _285_ (.A(_089_),
    .B(_202_),
    .X(_203_));
 sky130_fd_sc_hd__xor2_1 _286_ (.A(_201_),
    .B(_203_),
    .X(_204_));
 sky130_fd_sc_hd__and2_1 _287_ (.A(_200_),
    .B(_204_),
    .X(_205_));
 sky130_fd_sc_hd__nor2_1 _288_ (.A(_200_),
    .B(_204_),
    .Y(_206_));
 sky130_fd_sc_hd__nand2_1 _289_ (.A(net3),
    .B(_121_),
    .Y(_207_));
 sky130_fd_sc_hd__or2_1 _290_ (.A(net3),
    .B(_121_),
    .X(_208_));
 sky130_fd_sc_hd__a21oi_1 _291_ (.A1(_207_),
    .A2(_208_),
    .B1(_111_),
    .Y(_209_));
 sky130_fd_sc_hd__a31o_1 _292_ (.A1(_111_),
    .A2(_207_),
    .A3(_208_),
    .B1(_190_),
    .X(_210_));
 sky130_fd_sc_hd__o32a_1 _293_ (.A1(_198_),
    .A2(_205_),
    .A3(_206_),
    .B1(_209_),
    .B2(_210_),
    .X(_211_));
 sky130_fd_sc_hd__nand2_2 _294_ (.A(_197_),
    .B(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__or2_1 _295_ (.A(_195_),
    .B(_152_),
    .X(_213_));
 sky130_fd_sc_hd__a21oi_1 _296_ (.A1(_195_),
    .A2(_152_),
    .B1(_190_),
    .Y(_214_));
 sky130_fd_sc_hd__a22o_1 _297_ (.A1(_191_),
    .A2(_200_),
    .B1(_213_),
    .B2(_214_),
    .X(_215_));
 sky130_fd_sc_hd__and2_1 _298_ (.A(net3),
    .B(_192_),
    .X(_216_));
 sky130_fd_sc_hd__nor2_1 _299_ (.A(net3),
    .B(_192_),
    .Y(_217_));
 sky130_fd_sc_hd__xnor2_1 _300_ (.A(_121_),
    .B(_195_),
    .Y(_218_));
 sky130_fd_sc_hd__nor2_1 _301_ (.A(_089_),
    .B(_218_),
    .Y(_219_));
 sky130_fd_sc_hd__a21o_1 _302_ (.A1(_089_),
    .A2(_218_),
    .B1(_172_),
    .X(_220_));
 sky130_fd_sc_hd__o32a_2 _303_ (.A1(_191_),
    .A2(_216_),
    .A3(_217_),
    .B1(_219_),
    .B2(_220_),
    .X(_221_));
 sky130_fd_sc_hd__nor2_2 _304_ (.A(_215_),
    .B(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__xnor2_4 _305_ (.A(_212_),
    .B(_222_),
    .Y(_223_));
 sky130_fd_sc_hd__xor2_1 _306_ (.A(_197_),
    .B(_211_),
    .X(_224_));
 sky130_fd_sc_hd__xor2_2 _307_ (.A(net3),
    .B(_194_),
    .X(_225_));
 sky130_fd_sc_hd__xor2_1 _308_ (.A(_202_),
    .B(_100_),
    .X(_226_));
 sky130_fd_sc_hd__xnor2_1 _309_ (.A(_132_),
    .B(_226_),
    .Y(_227_));
 sky130_fd_sc_hd__xnor2_1 _310_ (.A(_225_),
    .B(_227_),
    .Y(_228_));
 sky130_fd_sc_hd__xor2_1 _311_ (.A(_121_),
    .B(_100_),
    .X(_229_));
 sky130_fd_sc_hd__xor2_1 _312_ (.A(_203_),
    .B(_229_),
    .X(_230_));
 sky130_fd_sc_hd__or3b_1 _313_ (.A(net9),
    .B(_230_),
    .C_N(_218_),
    .X(_231_));
 sky130_fd_sc_hd__o21bai_1 _314_ (.A1(_190_),
    .A2(_230_),
    .B1_N(_218_),
    .Y(_232_));
 sky130_fd_sc_hd__or2_1 _315_ (.A(_172_),
    .B(_195_),
    .X(_233_));
 sky130_fd_sc_hd__o2111a_1 _316_ (.A1(_191_),
    .A2(_228_),
    .B1(_231_),
    .C1(_232_),
    .D1(_233_),
    .X(_234_));
 sky130_fd_sc_hd__xor2_1 _317_ (.A(_195_),
    .B(_111_),
    .X(_235_));
 sky130_fd_sc_hd__xnor2_1 _318_ (.A(_192_),
    .B(_121_),
    .Y(_236_));
 sky130_fd_sc_hd__xnor2_1 _319_ (.A(_152_),
    .B(_236_),
    .Y(_237_));
 sky130_fd_sc_hd__mux2_1 _320_ (.A0(_235_),
    .A1(_237_),
    .S(_190_),
    .X(_238_));
 sky130_fd_sc_hd__xnor2_1 _321_ (.A(_195_),
    .B(_199_),
    .Y(_239_));
 sky130_fd_sc_hd__nand2_1 _322_ (.A(_201_),
    .B(_226_),
    .Y(_240_));
 sky130_fd_sc_hd__o21a_1 _323_ (.A1(_201_),
    .A2(_226_),
    .B1(net9),
    .X(_241_));
 sky130_fd_sc_hd__a22o_1 _324_ (.A1(_172_),
    .A2(_239_),
    .B1(_240_),
    .B2(_241_),
    .X(_242_));
 sky130_fd_sc_hd__nor2_1 _325_ (.A(_238_),
    .B(_242_),
    .Y(_243_));
 sky130_fd_sc_hd__xnor2_1 _326_ (.A(_234_),
    .B(_243_),
    .Y(_244_));
 sky130_fd_sc_hd__xnor2_1 _327_ (.A(_224_),
    .B(_244_),
    .Y(_245_));
 sky130_fd_sc_hd__xnor2_1 _328_ (.A(_223_),
    .B(_245_),
    .Y(_246_));
 sky130_fd_sc_hd__buf_2 _329_ (.A(_190_),
    .X(_247_));
 sky130_fd_sc_hd__xor2_1 _330_ (.A(_195_),
    .B(_142_),
    .X(_248_));
 sky130_fd_sc_hd__nand2_1 _331_ (.A(_247_),
    .B(_204_),
    .Y(_249_));
 sky130_fd_sc_hd__o21a_1 _332_ (.A1(_247_),
    .A2(_248_),
    .B1(_249_),
    .X(_250_));
 sky130_fd_sc_hd__nor2_1 _333_ (.A(_247_),
    .B(_225_),
    .Y(_251_));
 sky130_fd_sc_hd__a21o_1 _334_ (.A1(_247_),
    .A2(_201_),
    .B1(_251_),
    .X(_252_));
 sky130_fd_sc_hd__nor2_1 _335_ (.A(_250_),
    .B(_252_),
    .Y(_253_));
 sky130_fd_sc_hd__xnor2_2 _336_ (.A(_212_),
    .B(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__xor2_1 _337_ (.A(_202_),
    .B(_132_),
    .X(_255_));
 sky130_fd_sc_hd__nor2_1 _338_ (.A(_255_),
    .B(_162_),
    .Y(_256_));
 sky130_fd_sc_hd__a21o_1 _339_ (.A1(_255_),
    .A2(_162_),
    .B1(_191_),
    .X(_257_));
 sky130_fd_sc_hd__xor2_4 _340_ (.A(_192_),
    .B(_202_),
    .X(_258_));
 sky130_fd_sc_hd__xor2_2 _341_ (.A(_132_),
    .B(_258_),
    .X(_259_));
 sky130_fd_sc_hd__xor2_1 _342_ (.A(_100_),
    .B(_259_),
    .X(_260_));
 sky130_fd_sc_hd__a2bb2o_1 _343_ (.A1_N(_256_),
    .A2_N(_257_),
    .B1(_247_),
    .B2(_260_),
    .X(_261_));
 sky130_fd_sc_hd__nor2_1 _344_ (.A(_198_),
    .B(_230_),
    .Y(_000_));
 sky130_fd_sc_hd__nor2_1 _345_ (.A(_247_),
    .B(_259_),
    .Y(_001_));
 sky130_fd_sc_hd__or3_1 _346_ (.A(_191_),
    .B(_195_),
    .C(_259_),
    .X(_002_));
 sky130_fd_sc_hd__o31a_1 _347_ (.A1(_196_),
    .A2(_000_),
    .A3(_001_),
    .B1(_002_),
    .X(_003_));
 sky130_fd_sc_hd__nand2_1 _348_ (.A(_261_),
    .B(_003_),
    .Y(_004_));
 sky130_fd_sc_hd__nand2_1 _349_ (.A(_198_),
    .B(_239_),
    .Y(_005_));
 sky130_fd_sc_hd__xor2_1 _350_ (.A(net6),
    .B(_193_),
    .X(_006_));
 sky130_fd_sc_hd__xnor2_1 _351_ (.A(_005_),
    .B(_006_),
    .Y(_007_));
 sky130_fd_sc_hd__and2_1 _352_ (.A(_111_),
    .B(_258_),
    .X(_008_));
 sky130_fd_sc_hd__o21ai_1 _353_ (.A1(_111_),
    .A2(_258_),
    .B1(_190_),
    .Y(_009_));
 sky130_fd_sc_hd__xor2_1 _354_ (.A(_194_),
    .B(_100_),
    .X(_010_));
 sky130_fd_sc_hd__o22a_1 _355_ (.A1(_008_),
    .A2(_009_),
    .B1(_010_),
    .B2(_190_),
    .X(_011_));
 sky130_fd_sc_hd__nand2_1 _356_ (.A(_011_),
    .B(_182_),
    .Y(_012_));
 sky130_fd_sc_hd__xor2_1 _357_ (.A(_007_),
    .B(_012_),
    .X(_013_));
 sky130_fd_sc_hd__xnor2_1 _358_ (.A(_004_),
    .B(_013_),
    .Y(_014_));
 sky130_fd_sc_hd__xnor2_2 _359_ (.A(_254_),
    .B(_014_),
    .Y(_015_));
 sky130_fd_sc_hd__xor2_1 _360_ (.A(_225_),
    .B(_248_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _361_ (.A0(_203_),
    .A1(_016_),
    .S(_198_),
    .X(_017_));
 sky130_fd_sc_hd__and2_1 _362_ (.A(_229_),
    .B(_258_),
    .X(_018_));
 sky130_fd_sc_hd__o21ai_1 _363_ (.A1(_229_),
    .A2(_258_),
    .B1(_190_),
    .Y(_019_));
 sky130_fd_sc_hd__o22a_1 _364_ (.A1(_191_),
    .A2(_259_),
    .B1(_018_),
    .B2(_019_),
    .X(_020_));
 sky130_fd_sc_hd__xnor2_1 _365_ (.A(_194_),
    .B(_152_),
    .Y(_021_));
 sky130_fd_sc_hd__nor2_1 _366_ (.A(_191_),
    .B(_202_),
    .Y(_022_));
 sky130_fd_sc_hd__a21oi_1 _367_ (.A1(_247_),
    .A2(_021_),
    .B1(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__nand2_1 _368_ (.A(_020_),
    .B(_023_),
    .Y(_024_));
 sky130_fd_sc_hd__xor2_1 _369_ (.A(_243_),
    .B(_024_),
    .X(_025_));
 sky130_fd_sc_hd__xor2_2 _370_ (.A(_017_),
    .B(_025_),
    .X(_026_));
 sky130_fd_sc_hd__xor2_1 _371_ (.A(_254_),
    .B(_026_),
    .X(_027_));
 sky130_fd_sc_hd__nand2_1 _372_ (.A(_015_),
    .B(_027_),
    .Y(_028_));
 sky130_fd_sc_hd__xnor2_1 _373_ (.A(_254_),
    .B(_026_),
    .Y(_029_));
 sky130_fd_sc_hd__xnor2_1 _374_ (.A(_089_),
    .B(_021_),
    .Y(_030_));
 sky130_fd_sc_hd__mux2_1 _375_ (.A0(_259_),
    .A1(_030_),
    .S(_198_),
    .X(_031_));
 sky130_fd_sc_hd__nand2_1 _376_ (.A(_191_),
    .B(_236_),
    .Y(_032_));
 sky130_fd_sc_hd__o21ai_1 _377_ (.A1(_191_),
    .A2(_227_),
    .B1(_032_),
    .Y(_033_));
 sky130_fd_sc_hd__mux2_1 _378_ (.A0(_193_),
    .A1(_132_),
    .S(_172_),
    .X(_034_));
 sky130_fd_sc_hd__xor2_2 _379_ (.A(_202_),
    .B(_034_),
    .X(_035_));
 sky130_fd_sc_hd__nand2_1 _380_ (.A(_033_),
    .B(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__xnor2_1 _381_ (.A(_012_),
    .B(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__xnor2_2 _382_ (.A(_031_),
    .B(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__xnor2_4 _383_ (.A(_223_),
    .B(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__or3b_1 _384_ (.A(_246_),
    .B(_029_),
    .C_N(_039_),
    .X(_040_));
 sky130_fd_sc_hd__a21boi_1 _385_ (.A1(_246_),
    .A2(_028_),
    .B1_N(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__nand2_2 _386_ (.A(_182_),
    .B(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__or2_1 _387_ (.A(_039_),
    .B(_029_),
    .X(_043_));
 sky130_fd_sc_hd__xor2_1 _388_ (.A(_223_),
    .B(_245_),
    .X(_044_));
 sky130_fd_sc_hd__a21o_1 _389_ (.A1(_044_),
    .A2(_039_),
    .B1(_027_),
    .X(_045_));
 sky130_fd_sc_hd__a21o_1 _390_ (.A1(_045_),
    .A2(_040_),
    .B1(_015_),
    .X(_046_));
 sky130_fd_sc_hd__and2_1 _391_ (.A(_044_),
    .B(_015_),
    .X(_047_));
 sky130_fd_sc_hd__nand2_1 _392_ (.A(_039_),
    .B(_029_),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(_015_),
    .Y(_049_));
 sky130_fd_sc_hd__a22o_2 _394_ (.A1(_047_),
    .A2(_048_),
    .B1(_045_),
    .B2(_049_),
    .X(_050_));
 sky130_fd_sc_hd__a21o_1 _395_ (.A1(_043_),
    .A2(_046_),
    .B1(_050_),
    .X(_051_));
 sky130_fd_sc_hd__nand3_2 _396_ (.A(_050_),
    .B(_043_),
    .C(_046_),
    .Y(_052_));
 sky130_fd_sc_hd__a21oi_1 _397_ (.A1(_044_),
    .A2(_015_),
    .B1(_027_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_1 _398_ (.A(_246_),
    .B(_039_),
    .Y(_054_));
 sky130_fd_sc_hd__xnor2_2 _399_ (.A(_053_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__a21oi_1 _400_ (.A1(_039_),
    .A2(_027_),
    .B1(_015_),
    .Y(_056_));
 sky130_fd_sc_hd__nand2_1 _401_ (.A(_246_),
    .B(_039_),
    .Y(_057_));
 sky130_fd_sc_hd__xnor2_2 _402_ (.A(_056_),
    .B(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__xnor2_2 _403_ (.A(_055_),
    .B(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__a21oi_2 _404_ (.A1(_051_),
    .A2(_052_),
    .B1(_059_),
    .Y(_060_));
 sky130_fd_sc_hd__and3_1 _405_ (.A(_051_),
    .B(_052_),
    .C(_059_),
    .X(_061_));
 sky130_fd_sc_hd__nand3_1 _406_ (.A(_197_),
    .B(_051_),
    .C(_052_),
    .Y(_062_));
 sky130_fd_sc_hd__o31ai_1 _407_ (.A1(_221_),
    .A2(_060_),
    .A3(_061_),
    .B1(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__or4_1 _408_ (.A(_221_),
    .B(_062_),
    .C(_060_),
    .D(_061_),
    .X(_064_));
 sky130_fd_sc_hd__and3_1 _409_ (.A(_042_),
    .B(_063_),
    .C(_064_),
    .X(_065_));
 sky130_fd_sc_hd__a21oi_1 _410_ (.A1(_063_),
    .A2(_064_),
    .B1(_042_),
    .Y(_066_));
 sky130_fd_sc_hd__or2_2 _411_ (.A(_065_),
    .B(_066_),
    .X(_067_));
 sky130_fd_sc_hd__nand2_4 _412_ (.A(_261_),
    .B(_050_),
    .Y(_068_));
 sky130_fd_sc_hd__nand2_2 _413_ (.A(_011_),
    .B(_041_),
    .Y(_069_));
 sky130_fd_sc_hd__and2_1 _414_ (.A(_033_),
    .B(_055_),
    .X(_070_));
 sky130_fd_sc_hd__clkbuf_2 _415_ (.A(_070_),
    .X(_071_));
 sky130_fd_sc_hd__xnor2_2 _416_ (.A(_069_),
    .B(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__xnor2_1 _417_ (.A(_068_),
    .B(_072_),
    .Y(_073_));
 sky130_fd_sc_hd__mux2_2 _418_ (.A0(_028_),
    .A1(_047_),
    .S(_039_),
    .X(_074_));
 sky130_fd_sc_hd__nor2_4 _419_ (.A(_238_),
    .B(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__and3_1 _420_ (.A(_023_),
    .B(_043_),
    .C(_046_),
    .X(_076_));
 sky130_fd_sc_hd__buf_2 _421_ (.A(_076_),
    .X(_077_));
 sky130_fd_sc_hd__xor2_4 _422_ (.A(_075_),
    .B(_077_),
    .X(_078_));
 sky130_fd_sc_hd__xnor2_1 _423_ (.A(_073_),
    .B(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__nand2_1 _424_ (.A(_067_),
    .B(_079_),
    .Y(_080_));
 sky130_fd_sc_hd__o21a_1 _425_ (.A1(_067_),
    .A2(_079_),
    .B1(_198_),
    .X(_081_));
 sky130_fd_sc_hd__nor2_2 _426_ (.A(_242_),
    .B(_074_),
    .Y(_082_));
 sky130_fd_sc_hd__nor2b_2 _427_ (.A(_252_),
    .B_N(_059_),
    .Y(_083_));
 sky130_fd_sc_hd__xor2_1 _428_ (.A(_082_),
    .B(_083_),
    .X(_084_));
 sky130_fd_sc_hd__nand3_2 _429_ (.A(_020_),
    .B(_043_),
    .C(_046_),
    .Y(_085_));
 sky130_fd_sc_hd__xnor2_1 _430_ (.A(_062_),
    .B(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__xnor2_1 _431_ (.A(_084_),
    .B(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__buf_2 _432_ (.A(_247_),
    .X(_088_));
 sky130_fd_sc_hd__a22o_1 _433_ (.A1(_080_),
    .A2(_081_),
    .B1(_087_),
    .B2(_088_),
    .X(net10));
 sky130_fd_sc_hd__nor3_2 _434_ (.A(_221_),
    .B(_060_),
    .C(_061_),
    .Y(_090_));
 sky130_fd_sc_hd__xor2_1 _435_ (.A(_042_),
    .B(_090_),
    .X(_091_));
 sky130_fd_sc_hd__and3_1 _436_ (.A(_224_),
    .B(_051_),
    .C(_052_),
    .X(_092_));
 sky130_fd_sc_hd__clkbuf_2 _437_ (.A(_092_),
    .X(_093_));
 sky130_fd_sc_hd__xnor2_2 _438_ (.A(_072_),
    .B(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__or3_2 _439_ (.A(_215_),
    .B(_060_),
    .C(_061_),
    .X(_095_));
 sky130_fd_sc_hd__nand2_4 _440_ (.A(_035_),
    .B(_055_),
    .Y(_096_));
 sky130_fd_sc_hd__xnor2_1 _441_ (.A(_095_),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__xnor2_2 _442_ (.A(_094_),
    .B(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__nand2_1 _443_ (.A(_091_),
    .B(_098_),
    .Y(_099_));
 sky130_fd_sc_hd__or2_1 _444_ (.A(_091_),
    .B(_098_),
    .X(_101_));
 sky130_fd_sc_hd__xor2_1 _445_ (.A(_068_),
    .B(_071_),
    .X(_102_));
 sky130_fd_sc_hd__nand2b_4 _446_ (.A_N(_250_),
    .B(_059_),
    .Y(_103_));
 sky130_fd_sc_hd__xnor2_4 _447_ (.A(_069_),
    .B(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__xnor2_2 _448_ (.A(_095_),
    .B(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__xnor2_1 _449_ (.A(_102_),
    .B(_105_),
    .Y(_106_));
 sky130_fd_sc_hd__nand2_1 _450_ (.A(_063_),
    .B(_064_),
    .Y(_107_));
 sky130_fd_sc_hd__xor2_2 _451_ (.A(_107_),
    .B(_096_),
    .X(_108_));
 sky130_fd_sc_hd__nand2_1 _452_ (.A(_106_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__o21a_1 _453_ (.A1(_106_),
    .A2(_108_),
    .B1(_198_),
    .X(_110_));
 sky130_fd_sc_hd__a32o_1 _454_ (.A1(_088_),
    .A2(_099_),
    .A3(_101_),
    .B1(_109_),
    .B2(_110_),
    .X(net11));
 sky130_fd_sc_hd__xor2_1 _455_ (.A(_090_),
    .B(_094_),
    .X(_112_));
 sky130_fd_sc_hd__xnor2_2 _456_ (.A(_103_),
    .B(_112_),
    .Y(_113_));
 sky130_fd_sc_hd__nand2_1 _457_ (.A(_231_),
    .B(_232_),
    .Y(_114_));
 sky130_fd_sc_hd__nor2_1 _458_ (.A(_114_),
    .B(_058_),
    .Y(_115_));
 sky130_fd_sc_hd__xnor2_1 _459_ (.A(_096_),
    .B(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__xnor2_1 _460_ (.A(_068_),
    .B(_075_),
    .Y(_117_));
 sky130_fd_sc_hd__xnor2_1 _461_ (.A(_116_),
    .B(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__or2_1 _462_ (.A(_113_),
    .B(_118_),
    .X(_119_));
 sky130_fd_sc_hd__nand2_1 _463_ (.A(_113_),
    .B(_118_),
    .Y(_120_));
 sky130_fd_sc_hd__and2_1 _464_ (.A(_003_),
    .B(_050_),
    .X(_122_));
 sky130_fd_sc_hd__xor2_1 _465_ (.A(_078_),
    .B(_122_),
    .X(_123_));
 sky130_fd_sc_hd__o21ai_1 _466_ (.A1(_247_),
    .A2(_228_),
    .B1(_233_),
    .Y(_124_));
 sky130_fd_sc_hd__or2_1 _467_ (.A(_124_),
    .B(_058_),
    .X(_125_));
 sky130_fd_sc_hd__buf_2 _468_ (.A(_125_),
    .X(_126_));
 sky130_fd_sc_hd__xor2_2 _469_ (.A(_096_),
    .B(_126_),
    .X(_127_));
 sky130_fd_sc_hd__xor2_1 _470_ (.A(_085_),
    .B(_127_),
    .X(_128_));
 sky130_fd_sc_hd__xnor2_1 _471_ (.A(_123_),
    .B(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__xnor2_1 _472_ (.A(_105_),
    .B(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__nand2_1 _473_ (.A(_067_),
    .B(_130_),
    .Y(_131_));
 sky130_fd_sc_hd__o21a_1 _474_ (.A1(_067_),
    .A2(_130_),
    .B1(_198_),
    .X(_133_));
 sky130_fd_sc_hd__a32o_1 _475_ (.A1(_088_),
    .A2(_119_),
    .A3(_120_),
    .B1(_131_),
    .B2(_133_),
    .X(net12));
 sky130_fd_sc_hd__xor2_2 _476_ (.A(_077_),
    .B(_126_),
    .X(_134_));
 sky130_fd_sc_hd__xnor2_2 _477_ (.A(_085_),
    .B(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__xnor2_1 _478_ (.A(_083_),
    .B(_117_),
    .Y(_136_));
 sky130_fd_sc_hd__xnor2_1 _479_ (.A(_135_),
    .B(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__or2_1 _480_ (.A(_098_),
    .B(_137_),
    .X(_138_));
 sky130_fd_sc_hd__nand2_1 _481_ (.A(_098_),
    .B(_137_),
    .Y(_139_));
 sky130_fd_sc_hd__xnor2_1 _482_ (.A(_068_),
    .B(_077_),
    .Y(_140_));
 sky130_fd_sc_hd__xnor2_1 _483_ (.A(_082_),
    .B(_115_),
    .Y(_141_));
 sky130_fd_sc_hd__xnor2_1 _484_ (.A(_140_),
    .B(_141_),
    .Y(_143_));
 sky130_fd_sc_hd__xnor2_1 _485_ (.A(_126_),
    .B(_143_),
    .Y(_144_));
 sky130_fd_sc_hd__or2_1 _486_ (.A(_108_),
    .B(_144_),
    .X(_145_));
 sky130_fd_sc_hd__a21oi_1 _487_ (.A1(_108_),
    .A2(_144_),
    .B1(_088_),
    .Y(_146_));
 sky130_fd_sc_hd__a32o_1 _488_ (.A1(_088_),
    .A2(_138_),
    .A3(_139_),
    .B1(_145_),
    .B2(_146_),
    .X(net13));
 sky130_fd_sc_hd__xnor2_1 _489_ (.A(_078_),
    .B(_113_),
    .Y(_147_));
 sky130_fd_sc_hd__xnor2_1 _490_ (.A(_075_),
    .B(_141_),
    .Y(_148_));
 sky130_fd_sc_hd__xor2_1 _491_ (.A(_127_),
    .B(_148_),
    .X(_149_));
 sky130_fd_sc_hd__or2_1 _492_ (.A(_067_),
    .B(_149_),
    .X(_150_));
 sky130_fd_sc_hd__a21oi_1 _493_ (.A1(_067_),
    .A2(_149_),
    .B1(_088_),
    .Y(_151_));
 sky130_fd_sc_hd__a22o_1 _494_ (.A1(_088_),
    .A2(_147_),
    .B1(_150_),
    .B2(_151_),
    .X(net14));
 sky130_fd_sc_hd__xnor2_1 _495_ (.A(_083_),
    .B(_093_),
    .Y(_153_));
 sky130_fd_sc_hd__xnor2_1 _496_ (.A(_104_),
    .B(_153_),
    .Y(_154_));
 sky130_fd_sc_hd__or2_1 _497_ (.A(_123_),
    .B(_154_),
    .X(_155_));
 sky130_fd_sc_hd__nand2_1 _498_ (.A(_123_),
    .B(_154_),
    .Y(_156_));
 sky130_fd_sc_hd__xor2_2 _499_ (.A(_042_),
    .B(_122_),
    .X(_157_));
 sky130_fd_sc_hd__xor2_1 _500_ (.A(_104_),
    .B(_157_),
    .X(_158_));
 sky130_fd_sc_hd__xnor2_1 _501_ (.A(_090_),
    .B(_158_),
    .Y(_159_));
 sky130_fd_sc_hd__xnor2_1 _502_ (.A(_093_),
    .B(_116_),
    .Y(_160_));
 sky130_fd_sc_hd__xnor2_1 _503_ (.A(_135_),
    .B(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__nand2_1 _504_ (.A(_159_),
    .B(_161_),
    .Y(_163_));
 sky130_fd_sc_hd__o21a_1 _505_ (.A1(_159_),
    .A2(_161_),
    .B1(_088_),
    .X(_164_));
 sky130_fd_sc_hd__a32o_1 _506_ (.A1(_198_),
    .A2(_155_),
    .A3(_156_),
    .B1(_163_),
    .B2(_164_),
    .X(net15));
 sky130_fd_sc_hd__and3_1 _507_ (.A(_211_),
    .B(_051_),
    .C(_052_),
    .X(_165_));
 sky130_fd_sc_hd__o31ai_2 _508_ (.A1(_215_),
    .A2(_060_),
    .A3(_061_),
    .B1(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__or4_1 _509_ (.A(_215_),
    .B(_060_),
    .C(_061_),
    .D(_165_),
    .X(_167_));
 sky130_fd_sc_hd__nand3_1 _510_ (.A(_126_),
    .B(_166_),
    .C(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__a21o_1 _511_ (.A1(_166_),
    .A2(_167_),
    .B1(_126_),
    .X(_169_));
 sky130_fd_sc_hd__nand3_1 _512_ (.A(_107_),
    .B(_168_),
    .C(_169_),
    .Y(_170_));
 sky130_fd_sc_hd__a21o_1 _513_ (.A1(_168_),
    .A2(_169_),
    .B1(_107_),
    .X(_171_));
 sky130_fd_sc_hd__nand3_1 _514_ (.A(_148_),
    .B(_170_),
    .C(_171_),
    .Y(_173_));
 sky130_fd_sc_hd__a21o_1 _515_ (.A1(_170_),
    .A2(_171_),
    .B1(_148_),
    .X(_174_));
 sky130_fd_sc_hd__xnor2_1 _516_ (.A(_084_),
    .B(_160_),
    .Y(_175_));
 sky130_fd_sc_hd__xnor2_1 _517_ (.A(_157_),
    .B(_175_),
    .Y(_176_));
 sky130_fd_sc_hd__xnor2_1 _518_ (.A(_071_),
    .B(_134_),
    .Y(_177_));
 sky130_fd_sc_hd__xnor2_1 _519_ (.A(_103_),
    .B(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__nand2_1 _520_ (.A(_176_),
    .B(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__o21a_1 _521_ (.A1(_176_),
    .A2(_178_),
    .B1(_247_),
    .X(_180_));
 sky130_fd_sc_hd__a32o_1 _522_ (.A1(_198_),
    .A2(_173_),
    .A3(_174_),
    .B1(_179_),
    .B2(_180_),
    .X(net16));
 sky130_fd_sc_hd__a21oi_1 _523_ (.A1(_166_),
    .A2(_167_),
    .B1(_082_),
    .Y(_181_));
 sky130_fd_sc_hd__and3_1 _524_ (.A(_082_),
    .B(_166_),
    .C(_167_),
    .X(_183_));
 sky130_fd_sc_hd__or4_1 _525_ (.A(_065_),
    .B(_066_),
    .C(_181_),
    .D(_183_),
    .X(_184_));
 sky130_fd_sc_hd__o22ai_1 _526_ (.A1(_065_),
    .A2(_066_),
    .B1(_181_),
    .B2(_183_),
    .Y(_185_));
 sky130_fd_sc_hd__a21oi_1 _527_ (.A1(_184_),
    .A2(_185_),
    .B1(_127_),
    .Y(_186_));
 sky130_fd_sc_hd__a31o_1 _528_ (.A1(_127_),
    .A2(_184_),
    .A3(_185_),
    .B1(_088_),
    .X(_187_));
 sky130_fd_sc_hd__xor2_1 _529_ (.A(_042_),
    .B(_068_),
    .X(_188_));
 sky130_fd_sc_hd__xnor2_1 _530_ (.A(_113_),
    .B(_188_),
    .Y(_189_));
 sky130_fd_sc_hd__a2bb2o_1 _531_ (.A1_N(_186_),
    .A2_N(_187_),
    .B1(_189_),
    .B2(_088_),
    .X(net17));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(U[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(U[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(U[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(U[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(U[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(U[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(U[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(U[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(dec),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(S[0]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(S[1]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(S[2]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(S[3]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(S[4]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(S[5]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(S[6]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(S[7]));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_162 ();
endmodule
